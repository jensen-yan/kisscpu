module our(output cnt);
	initial begin
	    $display("Hello World");
	    $finish;
	end
	assign cnt = 1;
endmodule
